module IP2(input wire CLK,
            input wire RSTL,
            input wire PURGE,
            input wire [13:0] WADDRI,
            input wire BANKI,
            input wire WCEBI,
            input wire [127:0] DI,
            output wire [15:0] RADDRX,
            output wire [15:0] RADDRW,
            output wire [15:0] WADDRX,
            output wire BANKX,
            output wire BANKW,
            output wire RCEBW,
            output wire RCEBX,
            output wire WCEBX,
            output wire REQW,
            output wire WBUF_PURGE,
            output wire WBUF_EN,
            output wire [5:0] WBUF_EN_CTRL,
            output wire WBUF_ALL_EN,
            output wire WBUF_SWITCH,
            output wire FC_WEIGHT_EN,
            output wire NL_EN,
            output wire SHIFT_MODE,
            output wire [1:0] NL_SEL,
            output wire MAC_EN,
            output wire RESULT_REQ,
            output wire [3:0] OLSB,
            output wire RESULT_PURGE,
            output wire OUTPUT_EN,
            output wire [5:0] OUTPUT_EN_CTRL,
            output wire I_COMPARE_EN,
            output wire I_COMPARE_MODE,
            output wire I_COMPARE_SWITCH,
            output wire O_COMPARE_EN,
            output wire O_COMPARE_MODE,
            output wire O_COMPARE_SWITCH,
            output wire CAL_MODE,
            output wire CONV_FC_MODE,
            output wire FEEDBACK_MODE,
            output wire CONF_EN,
            output wire I_COMPARE_REGEN,
            output wire RCEBX0);
    
    wire [127:0] QI;
    wire RCEBI;
    wire [13:0] RADDRI;

    SEQUENCER sequencer_0(
        .CLK(CLK),
        .RSTL(RSTL),
        .PURGE(PURGE),
        //MEM Control for I
        .QI(QI),
        .RADDRI(RADDRI),
        .RCEBI(RCEBI),
        //MEM ADDR for X,W
        .RADDRX(RADDRX),
        .RADDRW(RADDRW),
        .WADDRX(WADDRX),
        //CTRL pins
        .BANKX(BANKX),
        .BANKW(BANKW),
        .RCEBX(RCEBX),
        .WCEBX(WCEBX),
        .RCEBW(RCEBW),
        .REQW(REQW),
        .WBUF_PURGE(WBUF_PURGE),
        .WBUF_EN(WBUF_EN),
        .WBUF_EN_CTRL(WBUF_EN_CTRL),
        .WBUF_ALL_EN(WBUF_ALL_EN),
        .WBUF_SWITCH(WBUF_SWITCH),
        .FC_WEIGHT_EN(FC_WEIGHT_EN),
        .NL_EN(NL_EN),
        .SHIFT_MODE(SHIFT_MODE),
        .NL_SEL(NL_SEL),
        .MAC_EN(MAC_EN),
        .RESULT_REQ(RESULT_REQ),
        .OLSB(OLSB),
        .RESULT_PURGE(RESULT_PURGE),
        .OUTPUT_EN(OUTPUT_EN),
        .OUTPUT_EN_CTRL(OUTPUT_EN_CTRL),
        .I_COMPARE_EN(I_COMPARE_EN),
        .I_COMPARE_MODE(I_COMPARE_MODE),
        .I_COMPARE_SWITCH(I_COMPARE_SWITCH),
        .O_COMPARE_EN(O_COMPARE_EN),
        .O_COMPARE_MODE(O_COMPARE_MODE),
        .O_COMPARE_SWITCH(O_COMPARE_SWITCH),
        .CAL_MODE(CAL_MODE),
        .CONV_FC_MODE(CONV_FC_MODE),
        .FEEDBACK_MODE(FEEDBACK_MODE),
        .CONF_EN(CONF_EN),
        .I_COMPARE_REGEN(I_COMPARE_REGEN),
        .RCEBX0(RCEBX0)
    );
    
    MEMI memi_0(
        .CLK(CLK),
        .RA(RADDRI),
        .RCEB(RCEBI),
        .BANK(BANKI),
        .WA(WADDRI),
        .WCEB(WCEBI),
        .DW(DI),
        .QW(QI)
    );
    
endmodule
